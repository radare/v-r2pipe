module r2pipe
