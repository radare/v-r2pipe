module main
import r2pipe

fn main() {
	res := r2pipe.cmd("x")
	println("hello: " + res)
}
